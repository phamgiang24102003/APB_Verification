package apb_seq_lib_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;

	import apb_agent_pkg::*;

	`include "apb_base_seq.sv"
	`include "apb_rd_seq.sv"
	`include "apb_wr_seq.sv"
	`include "apb_err_rd_seq.sv"
	`include "apb_err_wr_seq.sv"
endpackage
