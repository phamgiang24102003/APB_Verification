package apb_env_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;

	import apb_agent_pkg::*;

	`include"apb_env_cfg.sv"
	`include "apb_scoreboard.sv"
	`include "apb_env.sv"
endpackage
