module slave2 (
    input        PCLK,
    input        PRESETn,
    input        PSEL,
    input        PENABLE,
    input        PWRITE,
    input  [7:0] PADDR,
    input  [7:0] PWDATA,
    output [7:0] PRDATA2,
    output reg   PREADY
);

    reg [7:0] reg_addr;
    reg [7:0] mem2 [0:63];

    assign PRDATA2 = mem2[reg_addr];

    always @(*) begin
        if (!PRESETn)
            PREADY = 0;
        else if (PSEL && !PENABLE && !PWRITE)
            PREADY = 0;
        else if (PSEL && PENABLE && !PWRITE) begin
            PREADY    = 1;
            reg_addr  = PADDR;
        end else if (PSEL && !PENABLE && PWRITE)
            PREADY = 0;
        else if (PSEL && PENABLE && PWRITE) begin
            PREADY         = 1;
            mem2[PADDR]    = PWDATA;
        end else
            PREADY = 0;
    end

endmodule
