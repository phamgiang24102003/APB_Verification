package apb_test_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;

	import apb_agent_pkg::*;
	import apb_env_pkg::*;
	import apb_seq_lib_pkg::*;

	`include "apb_base_test.sv"
	`include "apb_test.sv"
endpackage
